-------------------------------------------------------------------------------
--
-- Title       : C4U
-- Design      : C4UD
-- Author      : tudorcampan@gmail.com
-- Company     : Sistemul Lamborghini SRL
--
-------------------------------------------------------------------------------
--
-- File        : D:\Proiect\C4UD\C4UD\src\C4U.vhd
-- Generated   : Fri May 22 21:04:18 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {C4U} architecture {C4U}}



entity C4U is
end C4U;

--}} End of automatically maintained section

architecture C4U of C4U is
begin

	 -- enter your statements here --

end C4U;
